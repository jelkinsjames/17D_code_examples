// Julian James
// 10/23/2022
// E E 371
// Lab 2 Task 2

// Implements both the internal RAM and controls the HEX displays.
// INPUTS: 1-bit clk, reset, wr_en, 4-bits wr_data 5-bits Wr_addr,
// OUTPUTS: 7-bit addrHEX1, addrHEX2, writeHEX, readHEX.
module RAMSystem (clk, reset, wr_en, wr_addr, wr_data, wr_addrHEX1, wr_addrHEX0, 
						re_addrHEX1, re_addrHEX0, wr_dataHEX, re_dataHEX);
	input logic clk, reset, wr_en;
	input logic [4:0] wr_addr;
	input logic [3:0] wr_data;
	output logic [6:0] wr_addrHEX1, wr_addrHEX0, re_addrHEX1, re_addrHEX0, wr_dataHEX, re_dataHEX;
	
	
	// The address that will be read, generated by the addrScroller.
	logic [4:0] addr_read;
	
	// Used to slow down the address scroller.
	logic [31:0] div_clk;
	
	// Used to pass the data read off the ram to the display.
	logic [3:0] re_data;
	
	
	
	clock_divider divider (.clock(clk), .divided_clocks(div_clk));
	
	addr_scroller scroller (.clk(div_clk[4]), .reset, .out(addr_read));
	

	// Outside inputs passed to ram and ram outputs passed to display.
	
	ram32x4 ram (.clock(clk), .data(wr_data), .rdaddress(addr_read), .wraddress(wr_addr), .wren(wr_en), .q(re_data));

	RAMDisplay display (.clk, . reset, .wr_addr, .wr_data, .re_addr(addr_read), .re_data, 
							  .re_addrHEX1, .re_addrHEX0, .wr_addrHEX1, .wr_addrHEX0, .wr_dataHEX, .re_dataHEX);
	
endmodule


`timescale 1 ps / 1 ps
module RAMSystem_testbench();
	logic clk, reset, wr_en;
	logic [3:0] wr_data;
	logic [4:0] wr_addr;
	logic [6:0] addrHEX1, addrHEX0, wrHEX, reHEX;
	
	RAMSystem dut (.clk, .reset, .wr_en, .wr_addr, .wr_data, .addrHEX1, .addrHEX0, .wrHEX, .reHEX);

	//Sets up the clock for use in the simulation.
	
	parameter clock_period = 100;
	initial begin
		clk <= 0;
		forever #(clock_period / 2) clk <= ~clk;
	end
	
	//Tests function of module as well as edgecases.
	initial begin
		reset <= 1; @(posedge clk);
		reset <= 0; @(posedge clk);
		wr_addr <= 5'b00000; wr_data <= 4'b0000; wr_en <= 0; repeat (16) @(posedge clk); 
		// writing data to address
		wr_en <= 1; wr_addr <= 5'b00001; wr_data <= 4'b0001; repeat(2) @(posedge clk); //hex should read 0 then 1
		// trying to write data to address when write <= 0
		wr_en <= 0; wr_addr <= 5'b00010; wr_data <= 4'b1000; repeat(2) @(posedge clk);
		//reading our old data
		wr_addr <= 5'b00001; @(posedge clk); // hex should read 1
		//changing old data again
		wr_en <= 1; repeat(3) @(posedge clk);
		
		$stop;
		
	end
endmodule